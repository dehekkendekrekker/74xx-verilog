(* extract_order = 4 *)
module MOD_74x08_1 (
    input A1,
    input B1,
    output Y1);

assign Y1 = A1 & B1;

endmodule
