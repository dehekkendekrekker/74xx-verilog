// 74x08 - Quad input AND Gate. Gate 1
module MOD_74x08_1 (
    input A,
    input B,
    output Y);

assign Y = A & B;

endmodule
