// 74x04 - Hex inverter. Gate 1
module MOD_74x04_1 (
    input A,
    output Y);

assign Y = ~A;

endmodule
