// 74x08 - Quad input OR Gate. Gates 1,2,3 and 4
module MOD_74x32_1 (
    input A,
    input B,
    output Y);

assign Y = A | B;

endmodule