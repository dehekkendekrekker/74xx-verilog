// 74x08 - Quad input XOR Gate.
module MOD_74x86_1 (
    input A,
    input B,
    output Y);

assign Y = A ^ B;

endmodule
